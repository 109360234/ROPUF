`timescale 1ns / 1ps
module R1(EN,Y1
    );
input EN;
output Y1;
wire w1,w2,w3,w4,w5;
	nand #1(w1,Y1,EN);
	not #1(w2,w1);
	not #1(w3,w2);
	not #1(w4,w3);
	not #1(Y1,w4);

endmodule
